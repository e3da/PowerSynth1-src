* 2018-10-31 14:56:17
R1 1 gnd 2.0
R2 2 3 4.0
R3 2 gnd 8.0
V1 1 2 DC 0 AC 1.0
V2 3 gnd DC 0 AC 1.0
.ac lin 1 1000Hz 1000Hz
.option post=2
.probe 
.option GENK=0
.end
